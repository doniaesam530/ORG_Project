

library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.segm_mips_const_pkg.all;

entity INSTRUCTION_MEMORY is
	port(
			RESET		: in	STD_LOGIC;						
  			READ_ADDR	: in	STD_LOGIC_VECTOR (INST_SIZE-1 downto 0);	
  			INST		: out	STD_LOGIC_VECTOR (INST_SIZE-1 downto 0)		
	);
end INSTRUCTION_MEMORY;


architecture INSTRUCTION_MEMORY_ARC of INSTRUCTION_MEMORY is
   
begin

	process (READ_ADDR)
	begin

		case READ_ADDR is
			when "00000000000000000000000000000000" => 
				INST <= "00000001010000000010000000100000";
			when "00000000000000000000000000000100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000001000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000001100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000010000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000010100" => 
				INST <= "00000000100000000001100000100000";
			when "00000000000000000000000000011000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000011100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000100000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000100100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000101000" => 
				INST <= "00000000011000110010000000100000";
			when "00000000000000000000000000101100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000110000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000110100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000111000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000000111100" => 
				INST <= "00000000100010110010000000100010";
			when "00000000000000000000000001000000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001000100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001001000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001001100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001010000" => 
				INST <= "00000000100000000100000000101010";
			when "00000000000000000000000001010100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001011000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001011100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001100000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001100100" => 
				INST <= "00010001000000010000000000001000";
			when "00000000000000000000000001101000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001101100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001110000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000001110100" => 
				INST <= "00000001100001010110000000100101";
			when "00000000000000000000000001111000" => 
				INST <= "00010000000000000000000000000100";
			when "00000000000000000000000001111100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010000000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010000100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010001000" => 
				INST <= "00000000011000110010000000100000";
			when "00000000000000000000000010001100" => 
				INST <= "00000000110000010011000000100000";
			when "00000000000000000000000010010000" => 
				INST <= "00000000101001010010100000100000";
			when "00000000000000000000000010010100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010011000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010011100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010100000" => 
				INST <= "00000000110001110100000000101010";
			when "00000000000000000000000010100100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010101000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010101100" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010110000" => 
				INST <= "00000000000000000000000000100010";
			when "00000000000000000000000010110100" => 
				INST <= "00010001000000011111111111010111";
			when others => 
				INST <= "11111111111111111111111111111111";
		end case;

	end process;

	
end INSTRUCTION_MEMORY_ARC;
