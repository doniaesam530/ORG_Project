library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity DataMemory is
	 port(
		 MemRead : in STD_LOGIC;
		 MemWrite : in STD_LOGIC;
		 Address : in STD_LOGIC_VECTOR(31 downto 0);
		 WriteData : in STD_LOGIC_VECTOR(31 downto 0);
		 ReadData : out STD_LOGIC_VECTOR(31 downto 0)
	     );
end DataMemory;



architecture DataMemory of DataMemory is
type RAM_16_x_32 is array(0 to 15) of std_logic_vector(31 downto 0);
signal DM : RAM_16_x_32:=(
"00000000000000000000001000001110",	--assume starts at 4
"00000000000000000000000000000000",
"00000000000000000000000000111100",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000",
"00000000000000000000000000000000"
);
begin
	process(memRead,memWrite)
	begin 
		if(memWrite='1') then
			DM((to_integer(unsigned(Address)))-4)<= WriteData;
		end if;
		if(memRead='1') then
			ReadData<=DM((to_integer(unsigned(Address)))-4);
		end if;
	end process;
	

end DataMemory;
